// =======================================================================
// Module:      RV32I Register File
// Project:     Ripple-32
// Description: The register file contains 32 registers, each 32 bits wide. 
// =======================================================================

module reg_file (
    input wire        clk,        
    input wire        rst_n
    // TODO add i/o ports for register file read/write
    
  );


endmodule